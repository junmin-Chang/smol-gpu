module shader_core(
    input test_input,
    output test_output
    );

assign test_output = ~test_input;

endmodule
